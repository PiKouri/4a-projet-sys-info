`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:36:08 04/16/2021 
// Design Name: 
// Module Name:    Memoire_Instructions 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Memoire_Instructions(
    input [7:0] addr,
    input CLK,
    output [31:0] OUT
    );


endmodule
